[program:cron]
command=/usr/sbin/crond
